module SC_regCLEAN #() (
	//////////// OUTPUTS //////////
	SC_RegCLEAN_OutBUS_InLow,
	//////////// INPUTS //////////
	SC_INITREGPOINT_7,
	SC_INITREGPOINT_6,
	SC_INITREGPOINT_5,
	SC_INITREGPOINT_4,
	SC_INITREGPOINT_3,
	SC_INITREGPOINT_2,
	SC_INITREGPOINT_1,
	SC_INITREGPOINT_0,
	SC_INITREGBACKG_7,
	SC_INITREGBACKG_6,
   SC_INITREGBACKG_5,
	SC_INITREGBACKG_4,
	SC_INITREGBACKG_3,
	SC_INITREGBACKG_2,
	SC_INITREGBACKG_1,
	SC_INITREGBACKG_0

);	

//=======================================================
//  PORT declarations
//=======================================================
output	SC_RegCLEAN_OutBUS_InLow;
input	[7:0]SC_INITREGPOINT_7;
input	[7:0]SC_INITREGPOINT_6;
input	[7:0]SC_INITREGPOINT_5;
input	[7:0]SC_INITREGPOINT_4;
input	[7:0]SC_INITREGPOINT_3;
input	[7:0]SC_INITREGPOINT_2;
input	[7:0]SC_INITREGPOINT_1;
input	[7:0]SC_INITREGPOINT_0;
input	[7:0]SC_INITREGBACKG_7;
input	[7:0]SC_INITREGBACKG_6;
input [7:0]SC_INITREGBACKG_5;
input	[7:0]SC_INITREGBACKG_4;
input	[7:0]SC_INITREGBACKG_3;
input	[7:0]SC_INITREGBACKG_2;
input	[7:0]SC_INITREGBACKG_1;
input	[7:0]SC_INITREGBACKG_0;

//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
always @(*)
begin
	if (SC_INITREGPOINT_7 | SC_INITREGBACKG_7 != 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_6 | SC_INITREGBACKG_6 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_5 | SC_INITREGBACKG_5 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_4 | SC_INITREGBACKG_4 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_3 | SC_INITREGBACKG_3 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_2 | SC_INITREGBACKG_2 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_1 | SC_INITREGBACKG_1 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else if (SC_INITREGPOINT_0 | SC_INITREGBACKG_0 == 8'b00000000)
		SC_RegCLEAN_OutBUS_InLow = 0;
	else
		SC_RegCLEAN_OutBUS_InLow = 1;
end

end
endmodule
